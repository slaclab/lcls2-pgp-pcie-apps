-------------------------------------------------------------------------------
-- File       : AppMigPkg.vhd
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2013-05-06
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description:
-- Package file for AXI DMA Controller
-------------------------------------------------------------------------------
-- This file is part of 'SLAC Firmware Standard Library'.
-- It is subject to the license terms in the LICENSE.txt file found in the 
-- top-level directory of this distribution and at: 
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html. 
-- No part of 'SLAC Firmware Standard Library', including this file, 
-- may be copied, modified, propagated, or distributed except according to 
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;


library surf;
use surf.StdRtlPkg.all;
use surf.AxiPkg.all;
use surf.AxiDmaPkg.all;

package AppMigPkg is

   constant BLOCK_BASE_SIZE_C : integer := 21; -- 2**17 = 128kB
   constant BLOCK_INDEX_SIZE_C : integer := 30 - BLOCK_BASE_SIZE_C;
   
   type MigConfigType is record
     blockSize   : slv(3 downto 0);
     blocksPause : slv(BLOCK_INDEX_SIZE_C-1 downto 0);
     inhibit     : sl;
     wrTagIndex  : slv(3 downto 0);
     rdEnable    : sl;
     rdAddr      : slv(BLOCK_INDEX_SIZE_C-1 downto 0);
   end record;

   -- Initialization constants
   constant MIG_CONFIG_INIT_C : MigConfigType := ( 
     blockSize   => toSlv(4,4),  -- 2MB
     blocksPause => toSlv(64,BLOCK_INDEX_SIZE_C),
     inhibit     => '1',
     wrTagIndex  => (others=>'0'),
     rdEnable    => '0',
     rdAddr      => (others=>'0') );

   -- Array
   type MigConfigArray is array (natural range<>) of MigConfigType;


   type MigStatusType is record
      memReady   : sl;
      wrIndex          : slv(BLOCK_INDEX_SIZE_C-1 downto 0);
      wcIndex          : slv(BLOCK_INDEX_SIZE_C-1 downto 0);
      rdIndex          : slv(BLOCK_INDEX_SIZE_C-1 downto 0);
      blocksQueued     : slv(BLOCK_INDEX_SIZE_C-1 downto 0);
      blocksFree       : slv(BLOCK_INDEX_SIZE_C-1 downto 0);
      writeQueCnt      : slv(7 downto 0);
      wid              : slv(7 downto 0);
      wdest            : slv(7 downto 0);
      rid              : slv(7 downto 0);
      rdest            : slv(7 downto 0);
      wrTagWc          : slv(1 downto 0);
      wrDescRetId      : slv(3 downto 0);
      wrTransAddr      : slv(15 downto 0);
      rdData           : slv(AXI_WRITE_DMA_DESC_RET_SIZE_C-1 downto 0);
      dmaWrStatus      : slv(7 downto 0);
   end record;

   constant MIG_STATUS_INIT_C : MigStatusType := (
      memReady        => '0',
      wrIndex         => (others=>'0'),
      wcIndex         => (others=>'0'),
      rdIndex         => (others=>'0'),
      blocksQueued    => (others=>'0'),
      blocksFree      => (others=>'0'),
      writeQueCnt     => (others=>'0'),
      wid             => (others=>'0'),
      wdest           => (others=>'0'),
      rid             => (others=>'0'),
      rdest           => (others=>'0'),
      wrTagWc         => (others=>'0'),
      wrDescRetId     => (others=>'0'),
      wrTransAddr     => (others=>'0'),
      rdData          => (others=>'0'),
      dmaWrStatus     => (others=>'0'));

   constant MIG_STATUS_BITS_C : integer := 71+5*BLOCK_INDEX_SIZE_C+AXI_WRITE_DMA_DESC_RET_SIZE_C;
   -- Array
   type MigStatusArray is array (natural range<>) of MigStatusType;

   function toSlv      (status : MigStatusType) return slv;
   function toMigStatus(vector : slv) return MigStatusType;

   constant APP2MIG_AXI_CONFIG_C : AxiConfigType := (
     ADDR_WIDTH_C => 32,
     DATA_BYTES_C => 16,
     ID_BITS_C    => 2,
     LEN_BITS_C   => 6 );

end package AppMigPkg;

package body AppMigPkg is

  function toSlv   (status : MigStatusType) return slv is
    variable vector : slv(MIG_STATUS_BITS_C-1 downto 0);
    variable i      : integer;
  begin
    assignSlv(i, vector, status.memReady);
    assignSlv(i, vector, status.wrIndex);
    assignSlv(i, vector, status.wcIndex);
    assignSlv(i, vector, status.rdIndex);
    assignSlv(i, vector, status.blocksQueued);
    assignSlv(i, vector, status.blocksFree);
    assignSlv(i, vector, status.writeQueCnt);
    assignSlv(i, vector, status.wid);
    assignSlv(i, vector, status.wdest);
    assignSlv(i, vector, status.rid);
    assignSlv(i, vector, status.rdest);
    assignSlv(i, vector, status.wrTagWc);
    assignSlv(i, vector, status.wrDescRetId);
    assignSlv(i, vector, status.wrTransAddr);
    assignSlv(i, vector, status.rdData);
    assignSlv(i, vector, status.dmaWrStatus);
    return vector;
  end function;

  function toMigStatus(vector : slv) return MigStatusType is
    variable status : MigStatusType;
    variable i      : integer := 0;
  begin
    assignRecord(i, vector, status.memReady);
    assignRecord(i, vector, status.wrIndex);
    assignRecord(i, vector, status.wcIndex);
    assignRecord(i, vector, status.rdIndex);
    assignRecord(i, vector, status.blocksQueued);
    assignRecord(i, vector, status.blocksFree);
    assignRecord(i, vector, status.writeQueCnt);
    assignRecord(i, vector, status.wid);
    assignRecord(i, vector, status.wdest);
    assignRecord(i, vector, status.rid);
    assignRecord(i, vector, status.rdest);
    assignRecord(i, vector, status.wrTagWc);
    assignRecord(i, vector, status.wrDescRetId);
    assignRecord(i, vector, status.wrTransAddr);
    assignRecord(i, vector, status.rdData);
    assignRecord(i, vector, status.dmaWrStatus);
    return status;
  end function;

end package body;
